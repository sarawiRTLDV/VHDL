-- Package Declaration Section
package microaddr_types is
	
	type cmd_t is (NONE, INC, JMP, JNZ, CALL, RET, OPJMP);
	
	
end package microaddr_types;